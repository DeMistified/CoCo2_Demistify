library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"c0fdc287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49c0fdc2",
    18 => x"48d8e4c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"d5e4c287",
    25 => x"d1e4c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e9c187f7",
    29 => x"e4c287f1",
    30 => x"e4c24dd5",
    31 => x"ad744cd5",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"731e741e",
    65 => x"c11e721e",
    66 => x"87cf048b",
    67 => x"02114812",
    68 => x"df4c87c9",
    69 => x"88749c98",
    70 => x"2687ec02",
    71 => x"264b264a",
    72 => x"1e4f264c",
    73 => x"73814873",
    74 => x"87c502a9",
    75 => x"f6055312",
    76 => x"1e4f2687",
    77 => x"4a711e73",
    78 => x"494b66c8",
    79 => x"99718bc1",
    80 => x"1287cf02",
    81 => x"08d4ff48",
    82 => x"c1497378",
    83 => x"0599718b",
    84 => x"4b2687f1",
    85 => x"5e0e4f26",
    86 => x"710e5c5b",
    87 => x"4cd4ff4a",
    88 => x"494b66cc",
    89 => x"99718bc1",
    90 => x"c387ce02",
    91 => x"526c7cff",
    92 => x"8bc14973",
    93 => x"f2059971",
    94 => x"264c2687",
    95 => x"1e4f264b",
    96 => x"d4ff1e73",
    97 => x"7bffc34b",
    98 => x"ffc34a6b",
    99 => x"c8496b7b",
   100 => x"c3b17232",
   101 => x"4a6b7bff",
   102 => x"b27131c8",
   103 => x"6b7bffc3",
   104 => x"7232c849",
   105 => x"264871b1",
   106 => x"0e4f264b",
   107 => x"5d5c5b5e",
   108 => x"ff4d710e",
   109 => x"48754cd4",
   110 => x"7098ffc3",
   111 => x"d8e4c27c",
   112 => x"87c805bf",
   113 => x"c94866d0",
   114 => x"58a6d430",
   115 => x"d84966d0",
   116 => x"c3487129",
   117 => x"7c7098ff",
   118 => x"d04966d0",
   119 => x"c3487129",
   120 => x"7c7098ff",
   121 => x"c84966d0",
   122 => x"c3487129",
   123 => x"7c7098ff",
   124 => x"c34866d0",
   125 => x"7c7098ff",
   126 => x"29d04975",
   127 => x"ffc34871",
   128 => x"6c7c7098",
   129 => x"fff0c94b",
   130 => x"abffc34a",
   131 => x"4987cf05",
   132 => x"4b6c7c71",
   133 => x"c5028ac1",
   134 => x"02ab7187",
   135 => x"487387f2",
   136 => x"4c264d26",
   137 => x"4f264b26",
   138 => x"ff49c01e",
   139 => x"ffc348d4",
   140 => x"c381c178",
   141 => x"04a9b7c8",
   142 => x"4f2687f1",
   143 => x"5c5b5e0e",
   144 => x"ffc00e5d",
   145 => x"4df7c1f0",
   146 => x"c0c0c0c1",
   147 => x"ff4bc0c0",
   148 => x"f8c487d6",
   149 => x"1ec04cdf",
   150 => x"cefd4975",
   151 => x"c186c487",
   152 => x"e5c005a8",
   153 => x"48d4ff87",
   154 => x"7378ffc3",
   155 => x"f0e1c01e",
   156 => x"fc49e9c1",
   157 => x"86c487f5",
   158 => x"ca059870",
   159 => x"48d4ff87",
   160 => x"c178ffc3",
   161 => x"fe87cb48",
   162 => x"8cc187de",
   163 => x"87c6ff05",
   164 => x"4d2648c0",
   165 => x"4b264c26",
   166 => x"5e0e4f26",
   167 => x"c00e5c5b",
   168 => x"c1c1f0ff",
   169 => x"48d4ff4c",
   170 => x"cb78ffc3",
   171 => x"f6f749dc",
   172 => x"c04bd387",
   173 => x"fb49741e",
   174 => x"86c487f1",
   175 => x"ca059870",
   176 => x"48d4ff87",
   177 => x"c178ffc3",
   178 => x"fd87cb48",
   179 => x"8bc187da",
   180 => x"87dfff05",
   181 => x"4c2648c0",
   182 => x"4f264b26",
   183 => x"00444d43",
   184 => x"43484453",
   185 => x"69616620",
   186 => x"000a216c",
   187 => x"52524549",
   188 => x"00000000",
   189 => x"00495053",
   190 => x"74697257",
   191 => x"61662065",
   192 => x"64656c69",
   193 => x"5e0e000a",
   194 => x"0e5d5c5b",
   195 => x"ff4dffc3",
   196 => x"d3fc4bd4",
   197 => x"1eeac687",
   198 => x"c1f0e1c0",
   199 => x"cafa49c8",
   200 => x"c186c487",
   201 => x"87c802a8",
   202 => x"c087effd",
   203 => x"87e8c148",
   204 => x"7087ccf9",
   205 => x"ffffcf49",
   206 => x"a9eac699",
   207 => x"fd87c802",
   208 => x"48c087d8",
   209 => x"7587d1c1",
   210 => x"4cf1c07b",
   211 => x"7087edfb",
   212 => x"ecc00298",
   213 => x"c01ec087",
   214 => x"fac1f0ff",
   215 => x"87cbf949",
   216 => x"987086c4",
   217 => x"7587da05",
   218 => x"75496b7b",
   219 => x"757b757b",
   220 => x"c17b757b",
   221 => x"c40299c0",
   222 => x"db48c187",
   223 => x"d748c087",
   224 => x"05acc287",
   225 => x"e0cb87ca",
   226 => x"87dbf449",
   227 => x"87c848c0",
   228 => x"fe058cc1",
   229 => x"48c087f6",
   230 => x"4c264d26",
   231 => x"4f264b26",
   232 => x"5c5b5e0e",
   233 => x"d0ff0e5d",
   234 => x"d0e5c04d",
   235 => x"c24cc0c1",
   236 => x"c148d8e4",
   237 => x"49f4cb78",
   238 => x"c787ecf3",
   239 => x"f97dc24b",
   240 => x"7dc387e6",
   241 => x"49741ec0",
   242 => x"c487e0f7",
   243 => x"05a8c186",
   244 => x"c24b87c1",
   245 => x"87cb05ab",
   246 => x"f349eccb",
   247 => x"48c087c9",
   248 => x"c187f6c0",
   249 => x"d4ff058b",
   250 => x"87dafc87",
   251 => x"58dce4c2",
   252 => x"cd059870",
   253 => x"c01ec187",
   254 => x"d0c1f0ff",
   255 => x"87ebf649",
   256 => x"d4ff86c4",
   257 => x"78ffc348",
   258 => x"c287eec4",
   259 => x"c258e0e4",
   260 => x"48d4ff7d",
   261 => x"c178ffc3",
   262 => x"264d2648",
   263 => x"264b264c",
   264 => x"5b5e0e4f",
   265 => x"710e5d5c",
   266 => x"4cffc34d",
   267 => x"744bd4ff",
   268 => x"48d0ff7b",
   269 => x"7478c3c4",
   270 => x"c01e757b",
   271 => x"d8c1f0ff",
   272 => x"87e7f549",
   273 => x"987086c4",
   274 => x"cb87cb02",
   275 => x"d6f149f8",
   276 => x"c048c187",
   277 => x"7b7487ee",
   278 => x"c87bfec3",
   279 => x"66d41ec0",
   280 => x"87cff349",
   281 => x"7b7486c4",
   282 => x"7b747b74",
   283 => x"4ae0dad8",
   284 => x"056b7b74",
   285 => x"8ac187c5",
   286 => x"7487f505",
   287 => x"48d0ff7b",
   288 => x"48c078c2",
   289 => x"4c264d26",
   290 => x"4f264b26",
   291 => x"5c5b5e0e",
   292 => x"86fc0e5d",
   293 => x"d4ff4b71",
   294 => x"c57ec04c",
   295 => x"4adfcdee",
   296 => x"6c7cffc3",
   297 => x"a8fec348",
   298 => x"87f8c005",
   299 => x"9b734d74",
   300 => x"d487cc02",
   301 => x"49731e66",
   302 => x"c487dbf2",
   303 => x"ff87d486",
   304 => x"d1c448d0",
   305 => x"4a66d478",
   306 => x"c17dffc3",
   307 => x"87f8058a",
   308 => x"c35aa6d8",
   309 => x"737c7cff",
   310 => x"87c5059b",
   311 => x"d048d0ff",
   312 => x"7e4ac178",
   313 => x"fe058ac1",
   314 => x"486e87f6",
   315 => x"4d268efc",
   316 => x"4b264c26",
   317 => x"731e4f26",
   318 => x"c04a711e",
   319 => x"48d4ff4b",
   320 => x"ff78ffc3",
   321 => x"c3c448d0",
   322 => x"48d4ff78",
   323 => x"7278ffc3",
   324 => x"f0ffc01e",
   325 => x"f249d1c1",
   326 => x"86c487d1",
   327 => x"d2059870",
   328 => x"1ec0c887",
   329 => x"fd4966cc",
   330 => x"86c487e2",
   331 => x"d0ff4b70",
   332 => x"7378c248",
   333 => x"264b2648",
   334 => x"5b5e0e4f",
   335 => x"c00e5d5c",
   336 => x"f0ffc01e",
   337 => x"f149c9c1",
   338 => x"1ed287e1",
   339 => x"49e8e4c2",
   340 => x"c887f9fc",
   341 => x"c14cc086",
   342 => x"acb7d284",
   343 => x"c287f804",
   344 => x"bf97e8e4",
   345 => x"99c0c349",
   346 => x"05a9c0c1",
   347 => x"c287e7c0",
   348 => x"bf97efe4",
   349 => x"c231d049",
   350 => x"bf97f0e4",
   351 => x"7232c84a",
   352 => x"f1e4c2b1",
   353 => x"b14abf97",
   354 => x"ffcf4c71",
   355 => x"c19cffff",
   356 => x"c134ca84",
   357 => x"e4c287e7",
   358 => x"49bf97f1",
   359 => x"99c631c1",
   360 => x"97f2e4c2",
   361 => x"b7c74abf",
   362 => x"c2b1722a",
   363 => x"bf97ede4",
   364 => x"9dcf4d4a",
   365 => x"97eee4c2",
   366 => x"9ac34abf",
   367 => x"e4c232ca",
   368 => x"4bbf97ef",
   369 => x"b27333c2",
   370 => x"97f0e4c2",
   371 => x"c0c34bbf",
   372 => x"2bb7c69b",
   373 => x"81c2b273",
   374 => x"307148c1",
   375 => x"48c14970",
   376 => x"4d703075",
   377 => x"84c14c72",
   378 => x"c0c89471",
   379 => x"cc06adb7",
   380 => x"b734c187",
   381 => x"b7c0c82d",
   382 => x"f4ff01ad",
   383 => x"26487487",
   384 => x"264c264d",
   385 => x"0e4f264b",
   386 => x"5d5c5b5e",
   387 => x"c286fc0e",
   388 => x"c048d0ed",
   389 => x"c8e5c278",
   390 => x"fb49c01e",
   391 => x"86c487d8",
   392 => x"c5059870",
   393 => x"c948c087",
   394 => x"4dc087d2",
   395 => x"48ccf2c2",
   396 => x"e5c278c1",
   397 => x"e2c04afe",
   398 => x"4bc849d4",
   399 => x"7087e7ea",
   400 => x"87c60598",
   401 => x"48ccf2c2",
   402 => x"e6c278c0",
   403 => x"e2c04ada",
   404 => x"4bc849e0",
   405 => x"7087cfea",
   406 => x"87c60598",
   407 => x"48ccf2c2",
   408 => x"f2c278c0",
   409 => x"c002bfcc",
   410 => x"ecc287fd",
   411 => x"c24dbfce",
   412 => x"bf9fc6ed",
   413 => x"d6c5487e",
   414 => x"c705a8ea",
   415 => x"ceecc287",
   416 => x"87ce4dbf",
   417 => x"e9ca486e",
   418 => x"c502a8d5",
   419 => x"c748c087",
   420 => x"e5c287ea",
   421 => x"49751ec8",
   422 => x"c487dbf9",
   423 => x"05987086",
   424 => x"48c087c5",
   425 => x"c287d5c7",
   426 => x"c04adae6",
   427 => x"c849ece2",
   428 => x"87f2e84b",
   429 => x"c8059870",
   430 => x"d0edc287",
   431 => x"d878c148",
   432 => x"fee5c287",
   433 => x"f8e2c04a",
   434 => x"e84bc849",
   435 => x"987087d8",
   436 => x"87c5c002",
   437 => x"e3c648c0",
   438 => x"c6edc287",
   439 => x"c149bf97",
   440 => x"c005a9d5",
   441 => x"edc287cd",
   442 => x"49bf97c7",
   443 => x"02a9eac2",
   444 => x"c087c5c0",
   445 => x"87c4c648",
   446 => x"97c8e5c2",
   447 => x"c3487ebf",
   448 => x"c002a8e9",
   449 => x"486e87ce",
   450 => x"02a8ebc3",
   451 => x"c087c5c0",
   452 => x"87e8c548",
   453 => x"97d3e5c2",
   454 => x"059949bf",
   455 => x"c287ccc0",
   456 => x"bf97d4e5",
   457 => x"02a9c249",
   458 => x"c087c5c0",
   459 => x"87ccc548",
   460 => x"97d5e5c2",
   461 => x"edc248bf",
   462 => x"4c7058cc",
   463 => x"c288c148",
   464 => x"c258d0ed",
   465 => x"bf97d6e5",
   466 => x"c2817549",
   467 => x"bf97d7e5",
   468 => x"7232c84a",
   469 => x"f1c27ea1",
   470 => x"786e48e8",
   471 => x"97d8e5c2",
   472 => x"f2c248bf",
   473 => x"edc258c0",
   474 => x"c202bfd0",
   475 => x"e6c287d3",
   476 => x"e2c04ada",
   477 => x"4bc849c8",
   478 => x"7087ebe5",
   479 => x"c5c00298",
   480 => x"c348c087",
   481 => x"edc287f6",
   482 => x"c24cbfc8",
   483 => x"c25cfcf1",
   484 => x"bf97ede5",
   485 => x"c231c849",
   486 => x"bf97ece5",
   487 => x"c249a14a",
   488 => x"bf97eee5",
   489 => x"7232d04a",
   490 => x"e5c249a1",
   491 => x"4abf97ef",
   492 => x"a17232d8",
   493 => x"c4f2c249",
   494 => x"fcf1c259",
   495 => x"f1c291bf",
   496 => x"c281bfe8",
   497 => x"c259f0f1",
   498 => x"bf97f5e5",
   499 => x"c232c84a",
   500 => x"bf97f4e5",
   501 => x"c24aa24b",
   502 => x"bf97f6e5",
   503 => x"7333d04b",
   504 => x"e5c24aa2",
   505 => x"4bbf97f7",
   506 => x"33d89bcf",
   507 => x"c24aa273",
   508 => x"c25af4f1",
   509 => x"c292748a",
   510 => x"7248f4f1",
   511 => x"c7c178a1",
   512 => x"dae5c287",
   513 => x"c849bf97",
   514 => x"d9e5c231",
   515 => x"a14abf97",
   516 => x"c731c549",
   517 => x"29c981ff",
   518 => x"59fcf1c2",
   519 => x"97dfe5c2",
   520 => x"32c84abf",
   521 => x"97dee5c2",
   522 => x"4aa24bbf",
   523 => x"5ac4f2c2",
   524 => x"bffcf1c2",
   525 => x"c2826e92",
   526 => x"c25af8f1",
   527 => x"c048f0f1",
   528 => x"ecf1c278",
   529 => x"78a17248",
   530 => x"48c4f2c2",
   531 => x"bff0f1c2",
   532 => x"c8f2c278",
   533 => x"f4f1c248",
   534 => x"edc278bf",
   535 => x"c002bfd0",
   536 => x"487487c9",
   537 => x"7e7030c4",
   538 => x"c287c9c0",
   539 => x"48bff8f1",
   540 => x"7e7030c4",
   541 => x"48d4edc2",
   542 => x"48c1786e",
   543 => x"4d268efc",
   544 => x"4b264c26",
   545 => x"00004f26",
   546 => x"33544146",
   547 => x"20202032",
   548 => x"00000000",
   549 => x"31544146",
   550 => x"20202036",
   551 => x"00000000",
   552 => x"33544146",
   553 => x"20202032",
   554 => x"00000000",
   555 => x"33544146",
   556 => x"20202032",
   557 => x"00000000",
   558 => x"31544146",
   559 => x"20202036",
   560 => x"5b5e0e00",
   561 => x"710e5d5c",
   562 => x"d0edc24a",
   563 => x"87cb02bf",
   564 => x"2bc74b72",
   565 => x"ffc14d72",
   566 => x"7287c99d",
   567 => x"722bc84b",
   568 => x"9dffc34d",
   569 => x"bfe8f1c2",
   570 => x"ccfac083",
   571 => x"d902abbf",
   572 => x"d0fac087",
   573 => x"c8e5c25b",
   574 => x"ef49731e",
   575 => x"86c487f8",
   576 => x"c5059870",
   577 => x"c048c087",
   578 => x"edc287e6",
   579 => x"d202bfd0",
   580 => x"c4497587",
   581 => x"c8e5c291",
   582 => x"cf4c6981",
   583 => x"ffffffff",
   584 => x"7587cb9c",
   585 => x"c291c249",
   586 => x"9f81c8e5",
   587 => x"48744c69",
   588 => x"4c264d26",
   589 => x"4f264b26",
   590 => x"5c5b5e0e",
   591 => x"86f40e5d",
   592 => x"c459a6c8",
   593 => x"80c84866",
   594 => x"c0487e70",
   595 => x"49c11e78",
   596 => x"87fdcc49",
   597 => x"4c7086c4",
   598 => x"fcc0029c",
   599 => x"d8edc287",
   600 => x"4966dc4a",
   601 => x"87e3ddff",
   602 => x"c0029870",
   603 => x"4a7487eb",
   604 => x"cb4966dc",
   605 => x"c7deff4b",
   606 => x"02987087",
   607 => x"1ec087db",
   608 => x"c4029c74",
   609 => x"c24dc087",
   610 => x"754dc187",
   611 => x"87c1cc49",
   612 => x"4c7086c4",
   613 => x"c4ff059c",
   614 => x"029c7487",
   615 => x"dc87f4c1",
   616 => x"486e49a4",
   617 => x"a4da7869",
   618 => x"4d66c449",
   619 => x"699f85c4",
   620 => x"d0edc27d",
   621 => x"87d202bf",
   622 => x"9f49a4d4",
   623 => x"ffc04969",
   624 => x"487199ff",
   625 => x"7e7030d0",
   626 => x"7ec087c2",
   627 => x"6d48496e",
   628 => x"c47d7080",
   629 => x"78c04866",
   630 => x"cc4966c4",
   631 => x"c4796d81",
   632 => x"81d04966",
   633 => x"a6c879c0",
   634 => x"c878c048",
   635 => x"66c44c66",
   636 => x"7482d44a",
   637 => x"7291c849",
   638 => x"41c049a1",
   639 => x"84c1796d",
   640 => x"04acb7c6",
   641 => x"c487e7ff",
   642 => x"c4c14966",
   643 => x"c179c081",
   644 => x"c087c248",
   645 => x"268ef448",
   646 => x"264c264d",
   647 => x"0e4f264b",
   648 => x"5d5c5b5e",
   649 => x"d04c710e",
   650 => x"496c4d66",
   651 => x"c2b97585",
   652 => x"4abfcced",
   653 => x"9972baff",
   654 => x"c0029971",
   655 => x"a4c487e4",
   656 => x"f9496b4b",
   657 => x"7b7087fb",
   658 => x"bfc8edc2",
   659 => x"71816c49",
   660 => x"c2b9757c",
   661 => x"4abfcced",
   662 => x"9972baff",
   663 => x"ff059971",
   664 => x"7c7587dc",
   665 => x"4c264d26",
   666 => x"4f264b26",
   667 => x"711e731e",
   668 => x"ecf1c24b",
   669 => x"a3c449bf",
   670 => x"c24a6a4a",
   671 => x"c8edc28a",
   672 => x"a17292bf",
   673 => x"ccedc249",
   674 => x"9a6b4abf",
   675 => x"c049a172",
   676 => x"c859d0fa",
   677 => x"e9711e66",
   678 => x"86c487dc",
   679 => x"c4059870",
   680 => x"c248c087",
   681 => x"2648c187",
   682 => x"1e4f264b",
   683 => x"4b711e73",
   684 => x"bfecf1c2",
   685 => x"4aa3c449",
   686 => x"8ac24a6a",
   687 => x"bfc8edc2",
   688 => x"49a17292",
   689 => x"bfccedc2",
   690 => x"729a6b4a",
   691 => x"fac049a1",
   692 => x"66c859d0",
   693 => x"c8e5711e",
   694 => x"7086c487",
   695 => x"87c40598",
   696 => x"87c248c0",
   697 => x"4b2648c1",
   698 => x"5e0e4f26",
   699 => x"0e5d5c5b",
   700 => x"4b7186e4",
   701 => x"4866ecc0",
   702 => x"a6cc28c9",
   703 => x"ccedc258",
   704 => x"b9ff49bf",
   705 => x"66c84871",
   706 => x"58a6d498",
   707 => x"986b4871",
   708 => x"c458a6d0",
   709 => x"a6c47ea3",
   710 => x"78bf6e48",
   711 => x"cc4866d0",
   712 => x"c605a866",
   713 => x"7b66c887",
   714 => x"d487c6c3",
   715 => x"ffc148a6",
   716 => x"ffffffff",
   717 => x"ff80c478",
   718 => x"d44ac078",
   719 => x"49724da3",
   720 => x"a17591c8",
   721 => x"4c66d049",
   722 => x"b7c08c69",
   723 => x"87cd04ac",
   724 => x"acb766d4",
   725 => x"dc87c603",
   726 => x"a6d85aa6",
   727 => x"c682c15c",
   728 => x"ff04aab7",
   729 => x"66d887d5",
   730 => x"a8b7c048",
   731 => x"d887d004",
   732 => x"91c84966",
   733 => x"2149a175",
   734 => x"69486e7b",
   735 => x"c087c978",
   736 => x"49a3cc7b",
   737 => x"7869486e",
   738 => x"6b4866c8",
   739 => x"58a6cc88",
   740 => x"bfc8edc2",
   741 => x"7090c848",
   742 => x"4866c87e",
   743 => x"c901a86e",
   744 => x"4866c887",
   745 => x"c003a86e",
   746 => x"c4c187fd",
   747 => x"bf6e7ea3",
   748 => x"7591c849",
   749 => x"66cc49a1",
   750 => x"49bf6e79",
   751 => x"a17591c8",
   752 => x"6681c449",
   753 => x"48a6d079",
   754 => x"d078bf6e",
   755 => x"a8c54866",
   756 => x"c487c705",
   757 => x"78c048a6",
   758 => x"66d087c8",
   759 => x"c880c148",
   760 => x"486e58a6",
   761 => x"c87866c4",
   762 => x"49731e66",
   763 => x"c487f0f8",
   764 => x"c8e5c286",
   765 => x"f949731e",
   766 => x"a3d087f2",
   767 => x"66f0c049",
   768 => x"268ee079",
   769 => x"264c264d",
   770 => x"0e4f264b",
   771 => x"0e5c5b5e",
   772 => x"4bc04a71",
   773 => x"c0029a72",
   774 => x"a2da87e0",
   775 => x"4b699f49",
   776 => x"bfd0edc2",
   777 => x"d487cf02",
   778 => x"699f49a2",
   779 => x"ffc04c49",
   780 => x"34d09cff",
   781 => x"4cc087c2",
   782 => x"9b73b374",
   783 => x"4a87df02",
   784 => x"edc28ac2",
   785 => x"9249bfc8",
   786 => x"bfecf1c2",
   787 => x"c2807248",
   788 => x"7158ccf2",
   789 => x"c230c448",
   790 => x"c058d8ed",
   791 => x"f1c287e9",
   792 => x"c24bbff0",
   793 => x"c248c8f2",
   794 => x"78bff4f1",
   795 => x"bfd0edc2",
   796 => x"c287c902",
   797 => x"49bfc8ed",
   798 => x"87c731c4",
   799 => x"bff8f1c2",
   800 => x"c231c449",
   801 => x"c259d8ed",
   802 => x"265bc8f2",
   803 => x"264b264c",
   804 => x"5b5e0e4f",
   805 => x"f00e5d5c",
   806 => x"59a6c886",
   807 => x"ffffffcf",
   808 => x"7ec04cf8",
   809 => x"d80266c4",
   810 => x"c4e5c287",
   811 => x"c278c048",
   812 => x"c248fce4",
   813 => x"78bfc8f2",
   814 => x"48c0e5c2",
   815 => x"bfc4f2c2",
   816 => x"e5edc278",
   817 => x"c250c048",
   818 => x"49bfd4ed",
   819 => x"bfc4e5c2",
   820 => x"03aa714a",
   821 => x"7287ccc4",
   822 => x"0599cf49",
   823 => x"c087eac0",
   824 => x"c248ccfa",
   825 => x"78bffce4",
   826 => x"1ec8e5c2",
   827 => x"bffce4c2",
   828 => x"fce4c249",
   829 => x"78a1c148",
   830 => x"f9dfff71",
   831 => x"c086c487",
   832 => x"c248c8fa",
   833 => x"cc78c8e5",
   834 => x"c8fac087",
   835 => x"e0c048bf",
   836 => x"ccfac080",
   837 => x"c4e5c258",
   838 => x"80c148bf",
   839 => x"58c8e5c2",
   840 => x"000e8827",
   841 => x"bf97bf00",
   842 => x"c2029d4d",
   843 => x"e5c387e5",
   844 => x"dec202ad",
   845 => x"c8fac087",
   846 => x"a3cb4bbf",
   847 => x"cf4c1149",
   848 => x"d2c105ac",
   849 => x"df497587",
   850 => x"cd89c199",
   851 => x"d8edc291",
   852 => x"4aa3c181",
   853 => x"a3c35112",
   854 => x"c551124a",
   855 => x"51124aa3",
   856 => x"124aa3c7",
   857 => x"4aa3c951",
   858 => x"a3ce5112",
   859 => x"d051124a",
   860 => x"51124aa3",
   861 => x"124aa3d2",
   862 => x"4aa3d451",
   863 => x"a3d65112",
   864 => x"d851124a",
   865 => x"51124aa3",
   866 => x"124aa3dc",
   867 => x"4aa3de51",
   868 => x"7ec15112",
   869 => x"7487fcc0",
   870 => x"0599c849",
   871 => x"7487edc0",
   872 => x"0599d049",
   873 => x"e0c087d3",
   874 => x"ccc00266",
   875 => x"c0497387",
   876 => x"700f66e0",
   877 => x"d3c00298",
   878 => x"c0056e87",
   879 => x"edc287c6",
   880 => x"50c048d8",
   881 => x"bfc8fac0",
   882 => x"87e9c248",
   883 => x"48e5edc2",
   884 => x"c27e50c0",
   885 => x"49bfd4ed",
   886 => x"bfc4e5c2",
   887 => x"04aa714a",
   888 => x"cf87f4fb",
   889 => x"f8ffffff",
   890 => x"c8f2c24c",
   891 => x"c8c005bf",
   892 => x"d0edc287",
   893 => x"fac102bf",
   894 => x"c0e5c287",
   895 => x"c0eb49bf",
   896 => x"c4e5c287",
   897 => x"48a6c458",
   898 => x"bfc0e5c2",
   899 => x"d0edc278",
   900 => x"dbc002bf",
   901 => x"4966c487",
   902 => x"a9749974",
   903 => x"87c8c002",
   904 => x"c048a6c8",
   905 => x"87e7c078",
   906 => x"c148a6c8",
   907 => x"87dfc078",
   908 => x"cf4966c4",
   909 => x"a999f8ff",
   910 => x"87c8c002",
   911 => x"c048a6cc",
   912 => x"87c5c078",
   913 => x"c148a6cc",
   914 => x"48a6c878",
   915 => x"c87866cc",
   916 => x"dec00566",
   917 => x"4966c487",
   918 => x"edc289c2",
   919 => x"c291bfc8",
   920 => x"48bfecf1",
   921 => x"e5c28071",
   922 => x"e5c258c0",
   923 => x"78c048c4",
   924 => x"c087d4f9",
   925 => x"ffffcf48",
   926 => x"f04cf8ff",
   927 => x"264d268e",
   928 => x"264b264c",
   929 => x"0000004f",
   930 => x"00000000",
   931 => x"ffffffff",
   932 => x"48d4ff1e",
   933 => x"6878ffc3",
   934 => x"1e4f2648",
   935 => x"c348d4ff",
   936 => x"d0ff78ff",
   937 => x"78e1c048",
   938 => x"d448d4ff",
   939 => x"1e4f2678",
   940 => x"c048d0ff",
   941 => x"4f2678e0",
   942 => x"87d4ff1e",
   943 => x"02994970",
   944 => x"fbc087c6",
   945 => x"87f105a9",
   946 => x"4f264871",
   947 => x"5c5b5e0e",
   948 => x"c04b710e",
   949 => x"87f8fe4c",
   950 => x"02994970",
   951 => x"c087f9c0",
   952 => x"c002a9ec",
   953 => x"fbc087f2",
   954 => x"ebc002a9",
   955 => x"b766cc87",
   956 => x"87c703ac",
   957 => x"c20266d0",
   958 => x"71537187",
   959 => x"87c20299",
   960 => x"cbfe84c1",
   961 => x"99497087",
   962 => x"c087cd02",
   963 => x"c702a9ec",
   964 => x"a9fbc087",
   965 => x"87d5ff05",
   966 => x"c30266d0",
   967 => x"7b97c087",
   968 => x"05a9ecc0",
   969 => x"4a7487c4",
   970 => x"4a7487c5",
   971 => x"728a0ac0",
   972 => x"264c2648",
   973 => x"1e4f264b",
   974 => x"7087d5fd",
   975 => x"a9f0c049",
   976 => x"c087c904",
   977 => x"c301a9f9",
   978 => x"89f0c087",
   979 => x"04a9c1c1",
   980 => x"dac187c9",
   981 => x"87c301a9",
   982 => x"7189f7c0",
   983 => x"0e4f2648",
   984 => x"5d5c5b5e",
   985 => x"7186f80e",
   986 => x"fc7ec04c",
   987 => x"4bc087ed",
   988 => x"97c0c0c1",
   989 => x"a9c049bf",
   990 => x"fc87cf04",
   991 => x"83c187fa",
   992 => x"97c0c0c1",
   993 => x"06ab49bf",
   994 => x"c0c187f1",
   995 => x"02bf97c0",
   996 => x"fbfb87cf",
   997 => x"99497087",
   998 => x"c087c602",
   999 => x"f105a9ec",
  1000 => x"fb4bc087",
  1001 => x"4d7087ea",
  1002 => x"c887e5fb",
  1003 => x"dffb58a6",
  1004 => x"c14a7087",
  1005 => x"49a4c883",
  1006 => x"ad496997",
  1007 => x"c987da05",
  1008 => x"699749a4",
  1009 => x"a966c449",
  1010 => x"ca87ce05",
  1011 => x"699749a4",
  1012 => x"c405aa49",
  1013 => x"d07ec187",
  1014 => x"adecc087",
  1015 => x"c087c602",
  1016 => x"c405adfb",
  1017 => x"c14bc087",
  1018 => x"fe026e7e",
  1019 => x"fefa87f5",
  1020 => x"f8487387",
  1021 => x"264d268e",
  1022 => x"264b264c",
  1023 => x"0000004f",
  1024 => x"1e731e00",
  1025 => x"c84bd4ff",
  1026 => x"d0ff4a66",
  1027 => x"78c5c848",
  1028 => x"c148d4ff",
  1029 => x"7b1178d4",
  1030 => x"f9058ac1",
  1031 => x"48d0ff87",
  1032 => x"4b2678c4",
  1033 => x"5e0e4f26",
  1034 => x"0e5d5c5b",
  1035 => x"7e7186f8",
  1036 => x"f2c21e6e",
  1037 => x"ffe349dc",
  1038 => x"7086c487",
  1039 => x"e4c40298",
  1040 => x"e8edc187",
  1041 => x"496e4cbf",
  1042 => x"c887d4fc",
  1043 => x"987058a6",
  1044 => x"c487c505",
  1045 => x"78c148a6",
  1046 => x"c548d0ff",
  1047 => x"48d4ff78",
  1048 => x"c478d5c1",
  1049 => x"89c14966",
  1050 => x"edc131c6",
  1051 => x"4abf97e0",
  1052 => x"ffb07148",
  1053 => x"ff7808d4",
  1054 => x"78c448d0",
  1055 => x"97d8f2c2",
  1056 => x"99d049bf",
  1057 => x"c587dd02",
  1058 => x"48d4ff78",
  1059 => x"c078d6c1",
  1060 => x"48d4ff4a",
  1061 => x"c178ffc3",
  1062 => x"aae0c082",
  1063 => x"ff87f204",
  1064 => x"78c448d0",
  1065 => x"c348d4ff",
  1066 => x"d0ff78ff",
  1067 => x"ff78c548",
  1068 => x"d3c148d4",
  1069 => x"ff78c178",
  1070 => x"78c448d0",
  1071 => x"06acb7c0",
  1072 => x"c287cbc2",
  1073 => x"4bbfe4f2",
  1074 => x"737e748c",
  1075 => x"ddc1029b",
  1076 => x"4dc0c887",
  1077 => x"abb7c08b",
  1078 => x"c887c603",
  1079 => x"c04da3c0",
  1080 => x"d8f2c24b",
  1081 => x"d049bf97",
  1082 => x"87cf0299",
  1083 => x"f2c21ec0",
  1084 => x"f7e549dc",
  1085 => x"7086c487",
  1086 => x"c287d84c",
  1087 => x"c21ec8e5",
  1088 => x"e549dcf2",
  1089 => x"4c7087e6",
  1090 => x"e5c21e75",
  1091 => x"f0fb49c8",
  1092 => x"7486c887",
  1093 => x"87c5059c",
  1094 => x"cac148c0",
  1095 => x"c21ec187",
  1096 => x"e349dcf2",
  1097 => x"86c487f9",
  1098 => x"fe059b73",
  1099 => x"4c6e87e3",
  1100 => x"06acb7c0",
  1101 => x"f2c287d1",
  1102 => x"78c048dc",
  1103 => x"78c080d0",
  1104 => x"f2c280f4",
  1105 => x"c078bfe8",
  1106 => x"fd01acb7",
  1107 => x"d0ff87f5",
  1108 => x"ff78c548",
  1109 => x"d3c148d4",
  1110 => x"ff78c078",
  1111 => x"78c448d0",
  1112 => x"c2c048c1",
  1113 => x"f848c087",
  1114 => x"264d268e",
  1115 => x"264b264c",
  1116 => x"5b5e0e4f",
  1117 => x"fc0e5d5c",
  1118 => x"c04d7186",
  1119 => x"04ad4c4b",
  1120 => x"c087e8c0",
  1121 => x"741edffd",
  1122 => x"87c4029c",
  1123 => x"87c24ac0",
  1124 => x"49724ac1",
  1125 => x"c487faeb",
  1126 => x"c17e7086",
  1127 => x"c2056e83",
  1128 => x"c14b7587",
  1129 => x"06ab7584",
  1130 => x"6e87d8ff",
  1131 => x"268efc48",
  1132 => x"264c264d",
  1133 => x"0e4f264b",
  1134 => x"0e5c5b5e",
  1135 => x"66cc4b71",
  1136 => x"4c87d802",
  1137 => x"028cf0c0",
  1138 => x"4a7487d8",
  1139 => x"d1028ac1",
  1140 => x"cd028a87",
  1141 => x"c9028a87",
  1142 => x"7387d987",
  1143 => x"87c6f949",
  1144 => x"1e7487d2",
  1145 => x"dac149c0",
  1146 => x"1e7487c2",
  1147 => x"d9c14973",
  1148 => x"86c887fa",
  1149 => x"4b264c26",
  1150 => x"5e0e4f26",
  1151 => x"0e5d5c5b",
  1152 => x"4c7186fc",
  1153 => x"c291de49",
  1154 => x"714dfcf3",
  1155 => x"026d9785",
  1156 => x"c287dcc1",
  1157 => x"49bfecf3",
  1158 => x"fd718174",
  1159 => x"7e7087d3",
  1160 => x"c0029848",
  1161 => x"f3c287f2",
  1162 => x"4a704bf0",
  1163 => x"fbfe49cb",
  1164 => x"4b7487f1",
  1165 => x"edc193cc",
  1166 => x"83c483ec",
  1167 => x"7bfcc9c1",
  1168 => x"c2c14974",
  1169 => x"7b7587fa",
  1170 => x"97e4edc1",
  1171 => x"c21e49bf",
  1172 => x"fd49f0f3",
  1173 => x"86c487e1",
  1174 => x"c2c14974",
  1175 => x"49c087e2",
  1176 => x"87fdc3c1",
  1177 => x"48d4f2c2",
  1178 => x"c04950c0",
  1179 => x"fc87c3e1",
  1180 => x"264d268e",
  1181 => x"264b264c",
  1182 => x"0000004f",
  1183 => x"64616f4c",
  1184 => x"2e676e69",
  1185 => x"00002e2e",
  1186 => x"61422080",
  1187 => x"00006b63",
  1188 => x"64616f4c",
  1189 => x"202e2a20",
  1190 => x"00000000",
  1191 => x"0000203a",
  1192 => x"61422080",
  1193 => x"00006b63",
  1194 => x"78452080",
  1195 => x"00007469",
  1196 => x"49204453",
  1197 => x"2e74696e",
  1198 => x"0000002e",
  1199 => x"00004b4f",
  1200 => x"544f4f42",
  1201 => x"20202020",
  1202 => x"004d4f52",
  1203 => x"711e731e",
  1204 => x"f3c2494b",
  1205 => x"7181bfec",
  1206 => x"7087d6fa",
  1207 => x"c4029a4a",
  1208 => x"e6e44987",
  1209 => x"ecf3c287",
  1210 => x"7378c048",
  1211 => x"87fac149",
  1212 => x"4f264b26",
  1213 => x"711e731e",
  1214 => x"4aa3c44b",
  1215 => x"87d0c102",
  1216 => x"dc028ac1",
  1217 => x"c0028a87",
  1218 => x"058a87f2",
  1219 => x"c287d3c1",
  1220 => x"02bfecf3",
  1221 => x"4887cbc1",
  1222 => x"f3c288c1",
  1223 => x"c1c158f0",
  1224 => x"ecf3c287",
  1225 => x"89c649bf",
  1226 => x"59f0f3c2",
  1227 => x"03a9b7c0",
  1228 => x"c287efc0",
  1229 => x"c048ecf3",
  1230 => x"87e6c078",
  1231 => x"bfe8f3c2",
  1232 => x"c287df02",
  1233 => x"48bfecf3",
  1234 => x"f3c280c1",
  1235 => x"87d258f0",
  1236 => x"bfe8f3c2",
  1237 => x"c287cb02",
  1238 => x"48bfecf3",
  1239 => x"f3c280c6",
  1240 => x"497358f0",
  1241 => x"4b2687c4",
  1242 => x"5e0e4f26",
  1243 => x"0e5d5c5b",
  1244 => x"a6d086f0",
  1245 => x"c8e5c259",
  1246 => x"c24cc04d",
  1247 => x"c148e8f3",
  1248 => x"48a6c878",
  1249 => x"7e7578c0",
  1250 => x"bfecf3c2",
  1251 => x"06a8c048",
  1252 => x"c887c0c1",
  1253 => x"7e755ca6",
  1254 => x"48c8e5c2",
  1255 => x"f2c00298",
  1256 => x"4d66c487",
  1257 => x"1edffdc0",
  1258 => x"c40266cc",
  1259 => x"c24cc087",
  1260 => x"744cc187",
  1261 => x"87d9e349",
  1262 => x"7e7086c4",
  1263 => x"66c885c1",
  1264 => x"cc80c148",
  1265 => x"f3c258a6",
  1266 => x"03adbfec",
  1267 => x"056e87c5",
  1268 => x"6e87d1ff",
  1269 => x"754cc04d",
  1270 => x"dcc3029d",
  1271 => x"dffdc087",
  1272 => x"0266cc1e",
  1273 => x"a6c887c7",
  1274 => x"c578c048",
  1275 => x"48a6c887",
  1276 => x"66c878c1",
  1277 => x"87d9e249",
  1278 => x"7e7086c4",
  1279 => x"c2029848",
  1280 => x"cb4987e4",
  1281 => x"49699781",
  1282 => x"c10299d0",
  1283 => x"497487d4",
  1284 => x"edc191cc",
  1285 => x"cbc181ec",
  1286 => x"81c879cc",
  1287 => x"7451ffc3",
  1288 => x"c291de49",
  1289 => x"714dfcf3",
  1290 => x"97c1c285",
  1291 => x"49a5c17d",
  1292 => x"c251e0c0",
  1293 => x"bf97d8ed",
  1294 => x"c187d202",
  1295 => x"4ba5c284",
  1296 => x"4ad8edc2",
  1297 => x"f3fe49db",
  1298 => x"d9c187d9",
  1299 => x"49a5cd87",
  1300 => x"84c151c0",
  1301 => x"6e4ba5c2",
  1302 => x"fe49cb4a",
  1303 => x"c187c4f3",
  1304 => x"497487c4",
  1305 => x"edc191cc",
  1306 => x"c7c181ec",
  1307 => x"edc279fa",
  1308 => x"02bf97d8",
  1309 => x"497487d8",
  1310 => x"84c191de",
  1311 => x"4bfcf3c2",
  1312 => x"edc28371",
  1313 => x"49dd4ad8",
  1314 => x"87d7f2fe",
  1315 => x"4b7487d8",
  1316 => x"f3c293de",
  1317 => x"a3cb83fc",
  1318 => x"c151c049",
  1319 => x"4a6e7384",
  1320 => x"f1fe49cb",
  1321 => x"66c887fd",
  1322 => x"cc80c148",
  1323 => x"acc758a6",
  1324 => x"87c5c003",
  1325 => x"e4fc056e",
  1326 => x"03acc787",
  1327 => x"c287e4c0",
  1328 => x"c048e8f3",
  1329 => x"cc497478",
  1330 => x"ecedc191",
  1331 => x"fac7c181",
  1332 => x"de497479",
  1333 => x"fcf3c291",
  1334 => x"c151c081",
  1335 => x"04acc784",
  1336 => x"c187dcff",
  1337 => x"c048c8ef",
  1338 => x"c180f750",
  1339 => x"c140d0d5",
  1340 => x"c878c8ca",
  1341 => x"f4cbc180",
  1342 => x"4966cc78",
  1343 => x"87c0f8c0",
  1344 => x"4d268ef0",
  1345 => x"4b264c26",
  1346 => x"731e4f26",
  1347 => x"494b711e",
  1348 => x"edc191cc",
  1349 => x"a1c881ec",
  1350 => x"e0edc14a",
  1351 => x"c9501248",
  1352 => x"c0c14aa1",
  1353 => x"501248c0",
  1354 => x"edc181ca",
  1355 => x"501148e4",
  1356 => x"97e4edc1",
  1357 => x"c01e49bf",
  1358 => x"87fbf149",
  1359 => x"e9f84973",
  1360 => x"268efc87",
  1361 => x"1e4f264b",
  1362 => x"f8c049c0",
  1363 => x"4f2687d3",
  1364 => x"494a711e",
  1365 => x"edc191cc",
  1366 => x"81c881ec",
  1367 => x"48d4f2c2",
  1368 => x"f0c05011",
  1369 => x"ecfe49a2",
  1370 => x"49c087e2",
  1371 => x"2687c3d5",
  1372 => x"d4ff1e4f",
  1373 => x"7affc34a",
  1374 => x"c048d0ff",
  1375 => x"7ade78e1",
  1376 => x"c8487a71",
  1377 => x"7a7028b7",
  1378 => x"b7d04871",
  1379 => x"717a7028",
  1380 => x"28b7d848",
  1381 => x"d0ff7a70",
  1382 => x"78e0c048",
  1383 => x"5e0e4f26",
  1384 => x"0e5d5c5b",
  1385 => x"4d7186f4",
  1386 => x"c191cc49",
  1387 => x"c881eced",
  1388 => x"a1ca4aa1",
  1389 => x"48a6c47e",
  1390 => x"bfd0f2c2",
  1391 => x"bf976e78",
  1392 => x"4c66c44b",
  1393 => x"48122c73",
  1394 => x"7058a6cc",
  1395 => x"c984c19c",
  1396 => x"49699781",
  1397 => x"c204acb7",
  1398 => x"6e4cc087",
  1399 => x"c84abf97",
  1400 => x"31724966",
  1401 => x"66c4b9ff",
  1402 => x"72487499",
  1403 => x"b14a7030",
  1404 => x"59d4f2c2",
  1405 => x"87f9fd71",
  1406 => x"f3c21ec7",
  1407 => x"c11ebfe4",
  1408 => x"c21eeced",
  1409 => x"bf97d4f2",
  1410 => x"87f4c149",
  1411 => x"f3c04975",
  1412 => x"8ee887ee",
  1413 => x"4c264d26",
  1414 => x"4f264b26",
  1415 => x"711e731e",
  1416 => x"f9fd494b",
  1417 => x"fd497387",
  1418 => x"4b2687f4",
  1419 => x"731e4f26",
  1420 => x"c24b711e",
  1421 => x"d6024aa3",
  1422 => x"058ac187",
  1423 => x"c287e2c0",
  1424 => x"02bfe4f3",
  1425 => x"c14887db",
  1426 => x"e8f3c288",
  1427 => x"c287d258",
  1428 => x"02bfe8f3",
  1429 => x"f3c287cb",
  1430 => x"c148bfe4",
  1431 => x"e8f3c280",
  1432 => x"c21ec758",
  1433 => x"1ebfe4f3",
  1434 => x"1eecedc1",
  1435 => x"97d4f2c2",
  1436 => x"87cc49bf",
  1437 => x"f2c04973",
  1438 => x"8ef487c6",
  1439 => x"4f264b26",
  1440 => x"5c5b5e0e",
  1441 => x"ccff0e5d",
  1442 => x"a6e8c086",
  1443 => x"48a6cc59",
  1444 => x"80c478c0",
  1445 => x"80c478c0",
  1446 => x"80c478c0",
  1447 => x"7866c8c1",
  1448 => x"78c180c4",
  1449 => x"78c180c4",
  1450 => x"48e8f3c2",
  1451 => x"dfff78c1",
  1452 => x"c3e087e9",
  1453 => x"d7dfff87",
  1454 => x"c04d7087",
  1455 => x"c102adfb",
  1456 => x"e4c087f3",
  1457 => x"e8c10566",
  1458 => x"66c4c187",
  1459 => x"6a82c44a",
  1460 => x"d0cac17e",
  1461 => x"20496e48",
  1462 => x"10412041",
  1463 => x"66c4c151",
  1464 => x"cad4c148",
  1465 => x"c7496a78",
  1466 => x"c1517581",
  1467 => x"c84966c4",
  1468 => x"dc51c181",
  1469 => x"78c248a6",
  1470 => x"4966c4c1",
  1471 => x"51c081c9",
  1472 => x"4966c4c1",
  1473 => x"51c081ca",
  1474 => x"1ed81ec1",
  1475 => x"81c8496a",
  1476 => x"87f8deff",
  1477 => x"c8c186c8",
  1478 => x"a8c04866",
  1479 => x"d487c701",
  1480 => x"78c148a6",
  1481 => x"c8c187cf",
  1482 => x"88c14866",
  1483 => x"c458a6dc",
  1484 => x"c3deff87",
  1485 => x"029d7587",
  1486 => x"d487f1cb",
  1487 => x"ccc14866",
  1488 => x"cb03a866",
  1489 => x"7ec087e6",
  1490 => x"87c4ddff",
  1491 => x"c1484d70",
  1492 => x"a6c888c6",
  1493 => x"02987058",
  1494 => x"4887d6c1",
  1495 => x"a6c888c9",
  1496 => x"02987058",
  1497 => x"4887d7c5",
  1498 => x"a6c888c1",
  1499 => x"02987058",
  1500 => x"4887f8c2",
  1501 => x"a6c888c3",
  1502 => x"02987058",
  1503 => x"c14887cf",
  1504 => x"58a6c888",
  1505 => x"c4029870",
  1506 => x"fec987f4",
  1507 => x"7ef0c087",
  1508 => x"87fcdbff",
  1509 => x"ecc04d70",
  1510 => x"87c202ad",
  1511 => x"ecc07e75",
  1512 => x"87cd02ad",
  1513 => x"87e8dbff",
  1514 => x"ecc04d70",
  1515 => x"f3ff05ad",
  1516 => x"66e4c087",
  1517 => x"87eac105",
  1518 => x"02adecc0",
  1519 => x"dbff87c4",
  1520 => x"1ec087ce",
  1521 => x"66dc1eca",
  1522 => x"c193cc4b",
  1523 => x"c48366cc",
  1524 => x"496c4ca3",
  1525 => x"87f4dbff",
  1526 => x"1ede1ec1",
  1527 => x"dbff496c",
  1528 => x"86d087ea",
  1529 => x"7bcad4c1",
  1530 => x"dc49a3c8",
  1531 => x"a3c95166",
  1532 => x"66e0c049",
  1533 => x"49a3ca51",
  1534 => x"66dc516e",
  1535 => x"c080c148",
  1536 => x"d458a6e0",
  1537 => x"66d84866",
  1538 => x"87cb04a8",
  1539 => x"c14866d4",
  1540 => x"58a6d880",
  1541 => x"d887fac7",
  1542 => x"88c14866",
  1543 => x"c758a6dc",
  1544 => x"daff87ef",
  1545 => x"4d7087d2",
  1546 => x"ff87e6c7",
  1547 => x"d087c8dc",
  1548 => x"66d058a6",
  1549 => x"87c606a8",
  1550 => x"cc48a6d0",
  1551 => x"dbff7866",
  1552 => x"ecc087f5",
  1553 => x"f5c105a8",
  1554 => x"66e4c087",
  1555 => x"87e5c105",
  1556 => x"cc4966d4",
  1557 => x"66c4c191",
  1558 => x"4aa1c481",
  1559 => x"a1c84c6a",
  1560 => x"5266cc4a",
  1561 => x"79d0d5c1",
  1562 => x"87e4d8ff",
  1563 => x"029d4d70",
  1564 => x"fbc087da",
  1565 => x"87d402ad",
  1566 => x"d8ff5475",
  1567 => x"4d7087d2",
  1568 => x"c7c0029d",
  1569 => x"adfbc087",
  1570 => x"87ecff05",
  1571 => x"c254e0c0",
  1572 => x"97c054c1",
  1573 => x"4866d47c",
  1574 => x"04a866d8",
  1575 => x"d487cbc0",
  1576 => x"80c14866",
  1577 => x"c558a6d8",
  1578 => x"66d887e7",
  1579 => x"dc88c148",
  1580 => x"dcc558a6",
  1581 => x"ffd7ff87",
  1582 => x"c54d7087",
  1583 => x"66cc87d3",
  1584 => x"66e4c048",
  1585 => x"f4c405a8",
  1586 => x"a6e8c087",
  1587 => x"ff78c048",
  1588 => x"7087e4d9",
  1589 => x"ded9ff7e",
  1590 => x"a6f0c087",
  1591 => x"a8ecc058",
  1592 => x"87c7c005",
  1593 => x"786e48a6",
  1594 => x"ff87c4c0",
  1595 => x"d487e1d6",
  1596 => x"91cc4966",
  1597 => x"4866c4c1",
  1598 => x"a6c88071",
  1599 => x"4a66c458",
  1600 => x"66c482c8",
  1601 => x"6e81ca49",
  1602 => x"66ecc051",
  1603 => x"6e81c149",
  1604 => x"7148c189",
  1605 => x"c1497030",
  1606 => x"7a977189",
  1607 => x"bfd0f2c2",
  1608 => x"97296e49",
  1609 => x"71484a6a",
  1610 => x"a6f4c098",
  1611 => x"4866c458",
  1612 => x"a6cc80c4",
  1613 => x"bf66c858",
  1614 => x"66e4c04c",
  1615 => x"a866cc48",
  1616 => x"87c5c002",
  1617 => x"c2c07ec0",
  1618 => x"6e7ec187",
  1619 => x"1ee0c01e",
  1620 => x"d5ff4974",
  1621 => x"86c887f6",
  1622 => x"b7c04d70",
  1623 => x"d4c106ad",
  1624 => x"c8847587",
  1625 => x"c049bf66",
  1626 => x"897481e0",
  1627 => x"dccac14b",
  1628 => x"defe714a",
  1629 => x"84c287ed",
  1630 => x"e8c07e74",
  1631 => x"80c14866",
  1632 => x"58a6ecc0",
  1633 => x"4966f0c0",
  1634 => x"a97081c1",
  1635 => x"87c5c002",
  1636 => x"c2c04cc0",
  1637 => x"744cc187",
  1638 => x"bf66cc1e",
  1639 => x"81e0c049",
  1640 => x"718966c4",
  1641 => x"4966c81e",
  1642 => x"87e0d4ff",
  1643 => x"b7c086c8",
  1644 => x"c5ff01a8",
  1645 => x"66e8c087",
  1646 => x"87d3c002",
  1647 => x"c94966c4",
  1648 => x"66e8c081",
  1649 => x"4866c451",
  1650 => x"78ded6c1",
  1651 => x"c487cec0",
  1652 => x"81c94966",
  1653 => x"66c451c2",
  1654 => x"dcd8c148",
  1655 => x"4866d478",
  1656 => x"04a866d8",
  1657 => x"d487cbc0",
  1658 => x"80c14866",
  1659 => x"c058a6d8",
  1660 => x"66d887d1",
  1661 => x"dc88c148",
  1662 => x"c6c058a6",
  1663 => x"f7d2ff87",
  1664 => x"cc4d7087",
  1665 => x"78c048a6",
  1666 => x"ff87c6c0",
  1667 => x"7087e9d2",
  1668 => x"66e0c04d",
  1669 => x"c080c148",
  1670 => x"7558a6e4",
  1671 => x"cbc0029d",
  1672 => x"4866d487",
  1673 => x"a866ccc1",
  1674 => x"87daf404",
  1675 => x"c74866d4",
  1676 => x"e1c003a8",
  1677 => x"4c66d487",
  1678 => x"48e8f3c2",
  1679 => x"497478c0",
  1680 => x"c4c191cc",
  1681 => x"a1c48166",
  1682 => x"c04a6a4a",
  1683 => x"84c17952",
  1684 => x"ff04acc7",
  1685 => x"e4c087e2",
  1686 => x"e2c00266",
  1687 => x"66c4c187",
  1688 => x"81d4c149",
  1689 => x"4a66c4c1",
  1690 => x"c082dcc1",
  1691 => x"d0d5c152",
  1692 => x"66c4c179",
  1693 => x"81d8c149",
  1694 => x"79e0cac1",
  1695 => x"c187d6c0",
  1696 => x"c14966c4",
  1697 => x"c4c181d4",
  1698 => x"d8c14a66",
  1699 => x"e8cac182",
  1700 => x"c7d5c17a",
  1701 => x"66c4c179",
  1702 => x"81e0c149",
  1703 => x"79eed8c1",
  1704 => x"87cbd0ff",
  1705 => x"ff4866d0",
  1706 => x"4d268ecc",
  1707 => x"4b264c26",
  1708 => x"c71e4f26",
  1709 => x"e4f3c21e",
  1710 => x"edc11ebf",
  1711 => x"f2c21eec",
  1712 => x"49bf97d4",
  1713 => x"c187f9ee",
  1714 => x"c049eced",
  1715 => x"f487ffe1",
  1716 => x"1e4f268e",
  1717 => x"48e0edc1",
  1718 => x"efc150c0",
  1719 => x"ff49bfd8",
  1720 => x"c087c3d5",
  1721 => x"1e4f2648",
  1722 => x"cdc71e73",
  1723 => x"f0f3c287",
  1724 => x"ff50c048",
  1725 => x"ffc348d4",
  1726 => x"f0cac178",
  1727 => x"e6d6fe49",
  1728 => x"dbe2fe87",
  1729 => x"02987087",
  1730 => x"ebfe87cd",
  1731 => x"987087f9",
  1732 => x"c187c402",
  1733 => x"c087c24a",
  1734 => x"029a724a",
  1735 => x"cac187c8",
  1736 => x"d6fe49fc",
  1737 => x"f3c287c1",
  1738 => x"78c048e4",
  1739 => x"48d4f2c2",
  1740 => x"fd4950c0",
  1741 => x"dafe87fc",
  1742 => x"9b4b7087",
  1743 => x"c187cf02",
  1744 => x"c75bc8ef",
  1745 => x"87f8de49",
  1746 => x"e0c049c1",
  1747 => x"f2c287d3",
  1748 => x"f4e1c087",
  1749 => x"dcf0c087",
  1750 => x"87f5ff87",
  1751 => x"4f264b26",
  1752 => x"00000000",
  1753 => x"00000000",
  1754 => x"00000001",
  1755 => x"000011fa",
  1756 => x"00002cfc",
  1757 => x"74000000",
  1758 => x"000011fa",
  1759 => x"00002d1a",
  1760 => x"74000000",
  1761 => x"000011fa",
  1762 => x"00002d38",
  1763 => x"74000000",
  1764 => x"000011fa",
  1765 => x"00002d56",
  1766 => x"74000000",
  1767 => x"000011fa",
  1768 => x"00002d74",
  1769 => x"74000000",
  1770 => x"000011fa",
  1771 => x"00002d92",
  1772 => x"74000000",
  1773 => x"000011fa",
  1774 => x"00002db0",
  1775 => x"74000000",
  1776 => x"00001550",
  1777 => x"00000000",
  1778 => x"74000000",
  1779 => x"000012f4",
  1780 => x"00000000",
  1781 => x"74000000",
  1782 => x"000012c0",
  1783 => x"db86fc1e",
  1784 => x"fc7e7087",
  1785 => x"1e4f268e",
  1786 => x"c048f0fe",
  1787 => x"7909cd78",
  1788 => x"1e4f2609",
  1789 => x"49dcefc1",
  1790 => x"4f2687ed",
  1791 => x"bff0fe1e",
  1792 => x"1e4f2648",
  1793 => x"c148f0fe",
  1794 => x"1e4f2678",
  1795 => x"c048f0fe",
  1796 => x"1e4f2678",
  1797 => x"52c04a71",
  1798 => x"0e4f2651",
  1799 => x"5d5c5b5e",
  1800 => x"7186f40e",
  1801 => x"7e6d974d",
  1802 => x"974ca5c1",
  1803 => x"a6c8486c",
  1804 => x"c4486e58",
  1805 => x"c505a866",
  1806 => x"c048ff87",
  1807 => x"caff87e6",
  1808 => x"49a5c287",
  1809 => x"714b6c97",
  1810 => x"6b974ba3",
  1811 => x"7e6c974b",
  1812 => x"80c1486e",
  1813 => x"c758a6c8",
  1814 => x"58a6cc98",
  1815 => x"fe7c9770",
  1816 => x"487387e1",
  1817 => x"4d268ef4",
  1818 => x"4b264c26",
  1819 => x"731e4f26",
  1820 => x"fe86f41e",
  1821 => x"bfe087d5",
  1822 => x"e0c0494b",
  1823 => x"c00299c0",
  1824 => x"4a7387ea",
  1825 => x"c29affc3",
  1826 => x"bf97e4f7",
  1827 => x"e6f7c249",
  1828 => x"c2517281",
  1829 => x"bf97e4f7",
  1830 => x"c1486e7e",
  1831 => x"58a6c880",
  1832 => x"a6cc98c7",
  1833 => x"e4f7c258",
  1834 => x"5066c848",
  1835 => x"7087cdfd",
  1836 => x"87cffd7e",
  1837 => x"4b268ef4",
  1838 => x"c21e4f26",
  1839 => x"fd49e4f7",
  1840 => x"f1c187d1",
  1841 => x"defc49ee",
  1842 => x"87e8c487",
  1843 => x"5e0e4f26",
  1844 => x"0e5d5c5b",
  1845 => x"7e7186fc",
  1846 => x"c24dd4ff",
  1847 => x"fc49e4f7",
  1848 => x"4b7087f9",
  1849 => x"04abb7c0",
  1850 => x"c387f5c2",
  1851 => x"c905abf0",
  1852 => x"ecf6c187",
  1853 => x"c278c148",
  1854 => x"e0c387d6",
  1855 => x"87c905ab",
  1856 => x"48f0f6c1",
  1857 => x"c7c278c1",
  1858 => x"f0f6c187",
  1859 => x"87c602bf",
  1860 => x"4ca3c0c2",
  1861 => x"4c7387c2",
  1862 => x"bfecf6c1",
  1863 => x"87e0c002",
  1864 => x"b7c44974",
  1865 => x"f6c19129",
  1866 => x"4a7481f4",
  1867 => x"92c29acf",
  1868 => x"307248c1",
  1869 => x"baff4a70",
  1870 => x"98694872",
  1871 => x"87db7970",
  1872 => x"b7c44974",
  1873 => x"f6c19129",
  1874 => x"4a7481f4",
  1875 => x"92c29acf",
  1876 => x"307248c3",
  1877 => x"69484a70",
  1878 => x"6e7970b0",
  1879 => x"87e4c005",
  1880 => x"c848d0ff",
  1881 => x"7dc578e1",
  1882 => x"bff0f6c1",
  1883 => x"c387c302",
  1884 => x"f6c17de0",
  1885 => x"c302bfec",
  1886 => x"7df0c387",
  1887 => x"d0ff7d73",
  1888 => x"78e0c048",
  1889 => x"48f0f6c1",
  1890 => x"f6c178c0",
  1891 => x"78c048ec",
  1892 => x"49e4f7c2",
  1893 => x"7087c4fa",
  1894 => x"abb7c04b",
  1895 => x"87cbfd03",
  1896 => x"8efc48c0",
  1897 => x"4c264d26",
  1898 => x"4f264b26",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"e4e4e4e4",
  1903 => x"e4e4e4e4",
  1904 => x"e4e4e4e4",
  1905 => x"e4e4e4e4",
  1906 => x"e4e4e4e4",
  1907 => x"e4e4e4e4",
  1908 => x"e4e4e4e4",
  1909 => x"e4e4e4e4",
  1910 => x"e4e4e4e4",
  1911 => x"e4e4e4e4",
  1912 => x"e4e4e4e4",
  1913 => x"e4e4e4e4",
  1914 => x"e4e4e4e4",
  1915 => x"e4e4e4e4",
  1916 => x"e4e4e4e4",
  1917 => x"724ac01e",
  1918 => x"c191c449",
  1919 => x"c081f4f6",
  1920 => x"d082c179",
  1921 => x"ee04aab7",
  1922 => x"0e4f2687",
  1923 => x"5d5c5b5e",
  1924 => x"f74d710e",
  1925 => x"4a7587f5",
  1926 => x"922ab7c4",
  1927 => x"82f4f6c1",
  1928 => x"9ccf4c75",
  1929 => x"496a94c2",
  1930 => x"c32b744b",
  1931 => x"7448c29b",
  1932 => x"ff4c7030",
  1933 => x"714874bc",
  1934 => x"f77a7098",
  1935 => x"487387c5",
  1936 => x"4c264d26",
  1937 => x"4f264b26",
  1938 => x"48d0ff1e",
  1939 => x"7178e1c8",
  1940 => x"08d4ff48",
  1941 => x"1e4f2678",
  1942 => x"c848d0ff",
  1943 => x"487178e1",
  1944 => x"7808d4ff",
  1945 => x"ff4866c4",
  1946 => x"267808d4",
  1947 => x"4a711e4f",
  1948 => x"1e4966c4",
  1949 => x"deff4972",
  1950 => x"48d0ff87",
  1951 => x"fc78e0c0",
  1952 => x"1e4f268e",
  1953 => x"4a711e73",
  1954 => x"abb7c24b",
  1955 => x"a387c803",
  1956 => x"ffc34a49",
  1957 => x"ce87c79a",
  1958 => x"c34a49a3",
  1959 => x"66c89aff",
  1960 => x"49721e49",
  1961 => x"fc87c6ff",
  1962 => x"264b268e",
  1963 => x"d0ff1e4f",
  1964 => x"78c9c848",
  1965 => x"d4ff4871",
  1966 => x"4f267808",
  1967 => x"494a711e",
  1968 => x"d0ff87eb",
  1969 => x"2678c848",
  1970 => x"1e731e4f",
  1971 => x"f7c24b71",
  1972 => x"c302bffc",
  1973 => x"87ebc287",
  1974 => x"c848d0ff",
  1975 => x"487378c9",
  1976 => x"ffb0e0c0",
  1977 => x"c27808d4",
  1978 => x"c048f0f7",
  1979 => x"0266c878",
  1980 => x"ffc387c5",
  1981 => x"c087c249",
  1982 => x"f8f7c249",
  1983 => x"0266cc59",
  1984 => x"d5c587c6",
  1985 => x"87c44ad5",
  1986 => x"4affffcf",
  1987 => x"5afcf7c2",
  1988 => x"48fcf7c2",
  1989 => x"4b2678c1",
  1990 => x"5e0e4f26",
  1991 => x"0e5d5c5b",
  1992 => x"f7c24d71",
  1993 => x"754bbff8",
  1994 => x"87cb029d",
  1995 => x"c191c849",
  1996 => x"714ac0fb",
  1997 => x"c187c482",
  1998 => x"c04ac0ff",
  1999 => x"7349124c",
  2000 => x"f4f7c299",
  2001 => x"b87148bf",
  2002 => x"7808d4ff",
  2003 => x"842bb7c1",
  2004 => x"04acb7c8",
  2005 => x"f7c287e7",
  2006 => x"c848bff0",
  2007 => x"f4f7c280",
  2008 => x"264d2658",
  2009 => x"264b264c",
  2010 => x"1e731e4f",
  2011 => x"4a134b71",
  2012 => x"87cb029a",
  2013 => x"e1fe4972",
  2014 => x"9a4a1387",
  2015 => x"2687f505",
  2016 => x"1e4f264b",
  2017 => x"bff0f7c2",
  2018 => x"f0f7c249",
  2019 => x"78a1c148",
  2020 => x"a9b7c0c4",
  2021 => x"ff87db03",
  2022 => x"f7c248d4",
  2023 => x"c278bff4",
  2024 => x"49bff0f7",
  2025 => x"48f0f7c2",
  2026 => x"c478a1c1",
  2027 => x"04a9b7c0",
  2028 => x"d0ff87e5",
  2029 => x"c278c848",
  2030 => x"c048fcf7",
  2031 => x"004f2678",
  2032 => x"00000000",
  2033 => x"00000000",
  2034 => x"5f000000",
  2035 => x"0000005f",
  2036 => x"00030300",
  2037 => x"00000303",
  2038 => x"147f7f14",
  2039 => x"00147f7f",
  2040 => x"6b2e2400",
  2041 => x"00123a6b",
  2042 => x"18366a4c",
  2043 => x"0032566c",
  2044 => x"594f7e30",
  2045 => x"40683a77",
  2046 => x"07040000",
  2047 => x"00000003",
  2048 => x"3e1c0000",
  2049 => x"00004163",
  2050 => x"63410000",
  2051 => x"00001c3e",
  2052 => x"1c3e2a08",
  2053 => x"082a3e1c",
  2054 => x"3e080800",
  2055 => x"0008083e",
  2056 => x"e0800000",
  2057 => x"00000060",
  2058 => x"08080800",
  2059 => x"00080808",
  2060 => x"60000000",
  2061 => x"00000060",
  2062 => x"18306040",
  2063 => x"0103060c",
  2064 => x"597f3e00",
  2065 => x"003e7f4d",
  2066 => x"7f060400",
  2067 => x"0000007f",
  2068 => x"71634200",
  2069 => x"00464f59",
  2070 => x"49632200",
  2071 => x"00367f49",
  2072 => x"13161c18",
  2073 => x"00107f7f",
  2074 => x"45672700",
  2075 => x"00397d45",
  2076 => x"4b7e3c00",
  2077 => x"00307949",
  2078 => x"71010100",
  2079 => x"00070f79",
  2080 => x"497f3600",
  2081 => x"00367f49",
  2082 => x"494f0600",
  2083 => x"001e3f69",
  2084 => x"66000000",
  2085 => x"00000066",
  2086 => x"e6800000",
  2087 => x"00000066",
  2088 => x"14080800",
  2089 => x"00222214",
  2090 => x"14141400",
  2091 => x"00141414",
  2092 => x"14222200",
  2093 => x"00080814",
  2094 => x"51030200",
  2095 => x"00060f59",
  2096 => x"5d417f3e",
  2097 => x"001e1f55",
  2098 => x"097f7e00",
  2099 => x"007e7f09",
  2100 => x"497f7f00",
  2101 => x"00367f49",
  2102 => x"633e1c00",
  2103 => x"00414141",
  2104 => x"417f7f00",
  2105 => x"001c3e63",
  2106 => x"497f7f00",
  2107 => x"00414149",
  2108 => x"097f7f00",
  2109 => x"00010109",
  2110 => x"417f3e00",
  2111 => x"007a7b49",
  2112 => x"087f7f00",
  2113 => x"007f7f08",
  2114 => x"7f410000",
  2115 => x"0000417f",
  2116 => x"40602000",
  2117 => x"003f7f40",
  2118 => x"1c087f7f",
  2119 => x"00416336",
  2120 => x"407f7f00",
  2121 => x"00404040",
  2122 => x"0c067f7f",
  2123 => x"007f7f06",
  2124 => x"0c067f7f",
  2125 => x"007f7f18",
  2126 => x"417f3e00",
  2127 => x"003e7f41",
  2128 => x"097f7f00",
  2129 => x"00060f09",
  2130 => x"61417f3e",
  2131 => x"00407e7f",
  2132 => x"097f7f00",
  2133 => x"00667f19",
  2134 => x"4d6f2600",
  2135 => x"00327b59",
  2136 => x"7f010100",
  2137 => x"0001017f",
  2138 => x"407f3f00",
  2139 => x"003f7f40",
  2140 => x"703f0f00",
  2141 => x"000f3f70",
  2142 => x"18307f7f",
  2143 => x"007f7f30",
  2144 => x"1c366341",
  2145 => x"4163361c",
  2146 => x"7c060301",
  2147 => x"0103067c",
  2148 => x"4d597161",
  2149 => x"00414347",
  2150 => x"7f7f0000",
  2151 => x"00004141",
  2152 => x"0c060301",
  2153 => x"40603018",
  2154 => x"41410000",
  2155 => x"00007f7f",
  2156 => x"03060c08",
  2157 => x"00080c06",
  2158 => x"80808080",
  2159 => x"00808080",
  2160 => x"03000000",
  2161 => x"00000407",
  2162 => x"54742000",
  2163 => x"00787c54",
  2164 => x"447f7f00",
  2165 => x"00387c44",
  2166 => x"447c3800",
  2167 => x"00004444",
  2168 => x"447c3800",
  2169 => x"007f7f44",
  2170 => x"547c3800",
  2171 => x"00185c54",
  2172 => x"7f7e0400",
  2173 => x"00000505",
  2174 => x"a4bc1800",
  2175 => x"007cfca4",
  2176 => x"047f7f00",
  2177 => x"00787c04",
  2178 => x"3d000000",
  2179 => x"0000407d",
  2180 => x"80808000",
  2181 => x"00007dfd",
  2182 => x"107f7f00",
  2183 => x"00446c38",
  2184 => x"3f000000",
  2185 => x"0000407f",
  2186 => x"180c7c7c",
  2187 => x"00787c0c",
  2188 => x"047c7c00",
  2189 => x"00787c04",
  2190 => x"447c3800",
  2191 => x"00387c44",
  2192 => x"24fcfc00",
  2193 => x"00183c24",
  2194 => x"243c1800",
  2195 => x"00fcfc24",
  2196 => x"047c7c00",
  2197 => x"00080c04",
  2198 => x"545c4800",
  2199 => x"00207454",
  2200 => x"7f3f0400",
  2201 => x"00004444",
  2202 => x"407c3c00",
  2203 => x"007c7c40",
  2204 => x"603c1c00",
  2205 => x"001c3c60",
  2206 => x"30607c3c",
  2207 => x"003c7c60",
  2208 => x"10386c44",
  2209 => x"00446c38",
  2210 => x"e0bc1c00",
  2211 => x"001c3c60",
  2212 => x"74644400",
  2213 => x"00444c5c",
  2214 => x"3e080800",
  2215 => x"00414177",
  2216 => x"7f000000",
  2217 => x"0000007f",
  2218 => x"77414100",
  2219 => x"0008083e",
  2220 => x"03010102",
  2221 => x"00010202",
  2222 => x"7f7f7f7f",
  2223 => x"007f7f7f",
  2224 => x"1c1c0808",
  2225 => x"7f7f3e3e",
  2226 => x"3e3e7f7f",
  2227 => x"08081c1c",
  2228 => x"7c181000",
  2229 => x"0010187c",
  2230 => x"7c301000",
  2231 => x"0010307c",
  2232 => x"60603010",
  2233 => x"00061e78",
  2234 => x"183c6642",
  2235 => x"0042663c",
  2236 => x"c26a3878",
  2237 => x"00386cc6",
  2238 => x"60000060",
  2239 => x"00600000",
  2240 => x"5c5b5e0e",
  2241 => x"86fc0e5d",
  2242 => x"f8c27e71",
  2243 => x"c04cbfc4",
  2244 => x"c41ec04b",
  2245 => x"c402ab66",
  2246 => x"c24dc087",
  2247 => x"754dc187",
  2248 => x"ee49731e",
  2249 => x"86c887e3",
  2250 => x"ef49e0c0",
  2251 => x"a4c487ec",
  2252 => x"f0496a4a",
  2253 => x"caf187f3",
  2254 => x"c184cc87",
  2255 => x"abb7c883",
  2256 => x"87cdff04",
  2257 => x"4d268efc",
  2258 => x"4b264c26",
  2259 => x"711e4f26",
  2260 => x"c8f8c24a",
  2261 => x"c8f8c25a",
  2262 => x"4978c748",
  2263 => x"2687e1fe",
  2264 => x"1e731e4f",
  2265 => x"b7c04a71",
  2266 => x"87d303aa",
  2267 => x"bfd8dbc2",
  2268 => x"c187c405",
  2269 => x"c087c24b",
  2270 => x"dcdbc24b",
  2271 => x"c287c45b",
  2272 => x"fc5adcdb",
  2273 => x"d8dbc248",
  2274 => x"c14a78bf",
  2275 => x"a2c0c19a",
  2276 => x"87e8ec49",
  2277 => x"4f264b26",
  2278 => x"c44a711e",
  2279 => x"49721e66",
  2280 => x"fc87e0eb",
  2281 => x"1e4f268e",
  2282 => x"c348d4ff",
  2283 => x"d0ff78ff",
  2284 => x"78e1c048",
  2285 => x"c148d4ff",
  2286 => x"c4487178",
  2287 => x"08d4ff30",
  2288 => x"48d0ff78",
  2289 => x"2678e0c0",
  2290 => x"5b5e0e4f",
  2291 => x"f40e5d5c",
  2292 => x"c87ec086",
  2293 => x"bfec48a6",
  2294 => x"c280fc78",
  2295 => x"78bfc4f8",
  2296 => x"bfccf8c2",
  2297 => x"4dbfe84c",
  2298 => x"bfd8dbc2",
  2299 => x"87dee349",
  2300 => x"d6e849c7",
  2301 => x"c2497087",
  2302 => x"87d00599",
  2303 => x"bfd0dbc2",
  2304 => x"c8b9ff49",
  2305 => x"99c19966",
  2306 => x"87fec102",
  2307 => x"cb49e8cf",
  2308 => x"4b7087ca",
  2309 => x"f2e749c7",
  2310 => x"05987087",
  2311 => x"66c887c9",
  2312 => x"0299c149",
  2313 => x"c887c3c1",
  2314 => x"bfec48a6",
  2315 => x"d8dbc278",
  2316 => x"d9e249bf",
  2317 => x"ca497387",
  2318 => x"987087ee",
  2319 => x"c287d702",
  2320 => x"49bfccdb",
  2321 => x"dbc2b9c1",
  2322 => x"fd7159d0",
  2323 => x"e8cf87d9",
  2324 => x"87c8ca49",
  2325 => x"49c74b70",
  2326 => x"7087f0e6",
  2327 => x"c6ff0598",
  2328 => x"4966c887",
  2329 => x"fe0599c1",
  2330 => x"dbc287fd",
  2331 => x"c14abfd8",
  2332 => x"dcdbc2ba",
  2333 => x"7a0afc5a",
  2334 => x"c19ac10a",
  2335 => x"e849a2c0",
  2336 => x"dac187fa",
  2337 => x"87c3e649",
  2338 => x"dbc27ec1",
  2339 => x"66c848d0",
  2340 => x"d8dbc278",
  2341 => x"e9c005bf",
  2342 => x"c3497587",
  2343 => x"1e7199ff",
  2344 => x"f3fb49c0",
  2345 => x"c8497587",
  2346 => x"1e7129b7",
  2347 => x"e7fb49c1",
  2348 => x"c386c887",
  2349 => x"d2e549fd",
  2350 => x"49fac387",
  2351 => x"c787cce5",
  2352 => x"497587fb",
  2353 => x"c899ffc3",
  2354 => x"b5712db7",
  2355 => x"c0029d75",
  2356 => x"a6c887e5",
  2357 => x"bfc8ff48",
  2358 => x"4966c878",
  2359 => x"bfd4dbc2",
  2360 => x"a9e0c289",
  2361 => x"87c5c003",
  2362 => x"d0c04dc0",
  2363 => x"d4dbc287",
  2364 => x"7866c848",
  2365 => x"c287c6c0",
  2366 => x"c048d4db",
  2367 => x"c8497578",
  2368 => x"cec00599",
  2369 => x"49f5c387",
  2370 => x"7087c0e4",
  2371 => x"0299c249",
  2372 => x"c287e4c0",
  2373 => x"02bfc8f8",
  2374 => x"4887cac0",
  2375 => x"f8c288c1",
  2376 => x"d0c058cc",
  2377 => x"4a66c487",
  2378 => x"6a82e0c1",
  2379 => x"87c5c002",
  2380 => x"7349ff4b",
  2381 => x"757ec10f",
  2382 => x"0599c449",
  2383 => x"c387cec0",
  2384 => x"c6e349f2",
  2385 => x"c2497087",
  2386 => x"edc00299",
  2387 => x"c8f8c287",
  2388 => x"c7487ebf",
  2389 => x"c003a8b7",
  2390 => x"486e87cb",
  2391 => x"f8c280c1",
  2392 => x"d3c058cc",
  2393 => x"4866c487",
  2394 => x"7080e0c1",
  2395 => x"02bf6e7e",
  2396 => x"4b87c5c0",
  2397 => x"0f7349fe",
  2398 => x"fdc37ec1",
  2399 => x"87cbe249",
  2400 => x"99c24970",
  2401 => x"87e6c002",
  2402 => x"bfc8f8c2",
  2403 => x"87c9c002",
  2404 => x"48c8f8c2",
  2405 => x"d3c078c0",
  2406 => x"4866c487",
  2407 => x"7080e0c1",
  2408 => x"02bf6e7e",
  2409 => x"4b87c5c0",
  2410 => x"0f7349fd",
  2411 => x"fac37ec1",
  2412 => x"87d7e149",
  2413 => x"99c24970",
  2414 => x"87eac002",
  2415 => x"bfc8f8c2",
  2416 => x"a8b7c748",
  2417 => x"87c9c003",
  2418 => x"48c8f8c2",
  2419 => x"d3c078c7",
  2420 => x"4866c487",
  2421 => x"7080e0c1",
  2422 => x"02bf6e7e",
  2423 => x"4b87c5c0",
  2424 => x"0f7349fc",
  2425 => x"48757ec1",
  2426 => x"cc98f0c3",
  2427 => x"987058a6",
  2428 => x"87cec005",
  2429 => x"e049dac1",
  2430 => x"497087d1",
  2431 => x"c10299c2",
  2432 => x"e8cf87ff",
  2433 => x"87d4c349",
  2434 => x"f8c24b70",
  2435 => x"50c048c0",
  2436 => x"97c0f8c2",
  2437 => x"d8c105bf",
  2438 => x"0566c887",
  2439 => x"c187cdc0",
  2440 => x"dfff49da",
  2441 => x"987087e5",
  2442 => x"87c5c102",
  2443 => x"494dbfe8",
  2444 => x"c899ffc3",
  2445 => x"b5712db7",
  2446 => x"bfd8dbc2",
  2447 => x"cddaff49",
  2448 => x"c2497387",
  2449 => x"987087e2",
  2450 => x"87c6c002",
  2451 => x"48c0f8c2",
  2452 => x"f8c250c1",
  2453 => x"05bf97c0",
  2454 => x"7587d6c0",
  2455 => x"99f0c349",
  2456 => x"87c8ff05",
  2457 => x"ff49dac1",
  2458 => x"7087e0de",
  2459 => x"fbfe0598",
  2460 => x"c8f8c287",
  2461 => x"cc4b49bf",
  2462 => x"8366c493",
  2463 => x"73714b6b",
  2464 => x"029c740f",
  2465 => x"6c87e9c0",
  2466 => x"87e4c002",
  2467 => x"ddff496c",
  2468 => x"497087f9",
  2469 => x"c00299c1",
  2470 => x"a4c487cb",
  2471 => x"c8f8c24b",
  2472 => x"4b6b49bf",
  2473 => x"0284c80f",
  2474 => x"6c87c5c0",
  2475 => x"87dcff05",
  2476 => x"c8c0026e",
  2477 => x"c8f8c287",
  2478 => x"c3f149bf",
  2479 => x"268ef487",
  2480 => x"264c264d",
  2481 => x"004f264b",
  2482 => x"00000010",
  2483 => x"00000000",
  2484 => x"00000000",
  2485 => x"00000000",
  2486 => x"00000000",
  2487 => x"ff4a711e",
  2488 => x"7249bfc8",
  2489 => x"4f2648a1",
  2490 => x"bfc8ff1e",
  2491 => x"c0c0fe89",
  2492 => x"a9c0c0c0",
  2493 => x"c087c401",
  2494 => x"c187c24a",
  2495 => x"2648724a",
  2496 => x"5b5e0e4f",
  2497 => x"710e5d5c",
  2498 => x"4cd4ff4b",
  2499 => x"c04866d0",
  2500 => x"ff49d678",
  2501 => x"c387f1dc",
  2502 => x"496c7cff",
  2503 => x"7199ffc3",
  2504 => x"f0c3494d",
  2505 => x"a9e0c199",
  2506 => x"c387cb05",
  2507 => x"486c7cff",
  2508 => x"66d098c3",
  2509 => x"ffc37808",
  2510 => x"494a6c7c",
  2511 => x"ffc331c8",
  2512 => x"714a6c7c",
  2513 => x"c84972b2",
  2514 => x"7cffc331",
  2515 => x"b2714a6c",
  2516 => x"31c84972",
  2517 => x"6c7cffc3",
  2518 => x"ffb2714a",
  2519 => x"e0c048d0",
  2520 => x"029b7378",
  2521 => x"7b7287c2",
  2522 => x"4d264875",
  2523 => x"4b264c26",
  2524 => x"261e4f26",
  2525 => x"5b5e0e4f",
  2526 => x"86f80e5c",
  2527 => x"a6c81e76",
  2528 => x"87fdfd49",
  2529 => x"4b7086c4",
  2530 => x"a8c4486e",
  2531 => x"87fbc203",
  2532 => x"f0c34a73",
  2533 => x"aad0c19a",
  2534 => x"c187c702",
  2535 => x"c205aae0",
  2536 => x"497387e9",
  2537 => x"c30299c8",
  2538 => x"87c6ff87",
  2539 => x"9cc34c73",
  2540 => x"c105acc2",
  2541 => x"66c487c4",
  2542 => x"7131c949",
  2543 => x"4a66c41e",
  2544 => x"c292ccc1",
  2545 => x"7249d0f8",
  2546 => x"ddccfe81",
  2547 => x"ff49d887",
  2548 => x"c887f5d9",
  2549 => x"e5c21ec0",
  2550 => x"e5fd49c8",
  2551 => x"d0ff87f8",
  2552 => x"78e0c048",
  2553 => x"1ec8e5c2",
  2554 => x"c14a66cc",
  2555 => x"f8c292cc",
  2556 => x"817249d0",
  2557 => x"87f3cafe",
  2558 => x"acc186cc",
  2559 => x"87cbc105",
  2560 => x"fd49eec0",
  2561 => x"c487c5e2",
  2562 => x"31c94966",
  2563 => x"66c41e71",
  2564 => x"92ccc14a",
  2565 => x"49d0f8c2",
  2566 => x"cbfe8172",
  2567 => x"e5c287cc",
  2568 => x"66c81ec8",
  2569 => x"92ccc14a",
  2570 => x"49d0f8c2",
  2571 => x"c8fe8172",
  2572 => x"49d787fa",
  2573 => x"87d0d8ff",
  2574 => x"c21ec0c8",
  2575 => x"fd49c8e5",
  2576 => x"cc87f0e3",
  2577 => x"48d0ff86",
  2578 => x"f878e0c0",
  2579 => x"264c268e",
  2580 => x"1e4f264b",
  2581 => x"b7c44a71",
  2582 => x"87ce03aa",
  2583 => x"ccc14972",
  2584 => x"d0f8c291",
  2585 => x"81c8c181",
  2586 => x"4f2679c0",
  2587 => x"5c5b5e0e",
  2588 => x"86fc0e5d",
  2589 => x"d4ff4a71",
  2590 => x"d44cc04b",
  2591 => x"b7c34d66",
  2592 => x"c2c201ad",
  2593 => x"029a7287",
  2594 => x"1e87ecc0",
  2595 => x"ccc14975",
  2596 => x"d0f8c291",
  2597 => x"c8807148",
  2598 => x"66c458a6",
  2599 => x"d7c2fe49",
  2600 => x"7086c487",
  2601 => x"87d40298",
  2602 => x"c8c1496e",
  2603 => x"6e79c181",
  2604 => x"6981c849",
  2605 => x"7587c54c",
  2606 => x"87d7fe49",
  2607 => x"c848d0ff",
  2608 => x"7bdd78e1",
  2609 => x"ffc34874",
  2610 => x"747b7098",
  2611 => x"29b7c849",
  2612 => x"ffc34871",
  2613 => x"747b7098",
  2614 => x"29b7d049",
  2615 => x"ffc34871",
  2616 => x"747b7098",
  2617 => x"28b7d848",
  2618 => x"7bc07b70",
  2619 => x"7b7b7b7b",
  2620 => x"7b7b7b7b",
  2621 => x"ff7b7b7b",
  2622 => x"e0c048d0",
  2623 => x"dc1e7578",
  2624 => x"e8d5ff49",
  2625 => x"fc86c487",
  2626 => x"264d268e",
  2627 => x"264b264c",
  2628 => x"001bf34f",
  2629 => x"001bf300",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
